`timescale 1ns/1ps
`default_nettype none

module inputqueue #(
    //params here
)(
// inputs/outputs declared here
);
//logic here
endmodule